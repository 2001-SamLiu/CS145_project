`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/04/07 08:14:41
// Design Name: 
// Module Name: dataMemory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dataMemory(
    input Clk,
    input [31:0] address,
    input [31:0] writeData,
    input memWrite,
    input memRead,
    output [31:0] readData
    );
    reg[31:0] memFile[0:63];
    integer i;
    initial begin
    for(i=0;i<64;i=i+1)
    memFile[i]=0;
    end
    reg[31:0] ReadData=0;
    assign readData=ReadData;
    always@(address)
    begin
    if(memRead==1)
    ReadData=memFile[address];
    end
    always@(negedge Clk)
    begin
    if(memWrite)
    memFile[address]=writeData;
    end
endmodule
